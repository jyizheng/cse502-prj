/* Instruction-Fetch */
module INF();

endmodule

/* vim: set ts=4 sw=0 tw=0 noet : */
