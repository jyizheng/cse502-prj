module Decoder ();
endmodule

