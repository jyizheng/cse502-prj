`ifndef _MEMORY_SVH_
`define _MEMORY_SVH_

`define MEM_TAG_I	8`h01
`define MEM_TAG_D	8`h04

`endif
