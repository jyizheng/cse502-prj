
`ifndef _CACHE_SVH_
`define _CACHE_SVH_ 1

`define CL_ACC_V	63
`define CL_ACC_D	62
`define CL_ACC_T	61	/* Timing bit for LRU */

`define CL_ACC_T_LSB	0
`define CL_ACC_T_MSB	48

`define CL_WEN_ALL	8'hFF

`endif
/* vim: set ts=4 sw=0 tw=0 noet : */
