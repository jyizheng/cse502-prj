`ifndef _GLOBAL_SVH_
`define _GLOBAL_SVH_ 1

`define GLB_REG_NUM	32

`endif

/* vim: set ts=4 sw=0 tw=0 noet : */
